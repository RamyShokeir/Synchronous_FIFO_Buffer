package  sync_fifo_pkg;

parameter  BUS_WIDTH = 32 ;
parameter  BUFFER_DEPTH = 256;

endpackage