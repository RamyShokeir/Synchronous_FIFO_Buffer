package  shared_pkg;

parameter  BUS_WIDTH = 32 ;
parameter  BUFFER_DEPTH = 16;
static int error_count;
static int correct_count;
bit test_finished;
endpackage